library verilog;
use verilog.vl_types.all;
entity dut_if is
    port(
        clk             : in     vl_logic;
        rst             : in     vl_logic
    );
end dut_if;
