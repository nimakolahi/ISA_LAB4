library verilog;
use verilog.vl_types.all;
entity DUT is
    port(
        state           : out    vl_logic
    );
end DUT;
